`timescale 1ps / 1ps
module tb_syn_arc4 ();


endmodule : tb_syn_arc4
