module tb_rtl_arc4();

`timescale 1ps / 1ps

endmodule: tb_rtl_arc4
