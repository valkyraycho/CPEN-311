`timescale 1ps / 1ps
module tb_rtl_prga();




endmodule: tb_rtl_prga
