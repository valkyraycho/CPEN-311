`timescale 1ps / 1ps
module tb_syn_prga ();


endmodule : tb_syn_prga
