module tb_syn_prga();

`timescale 1ps / 1ps

endmodule: tb_syn_prga
