module tb_syn_task3();

`timescale 1ps / 1ps

endmodule: tb_syn_task3
