module tb_syn_arc4();

`timescale 1ps / 1ps

endmodule: tb_syn_arc4
